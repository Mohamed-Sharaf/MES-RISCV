module fp_mv (
    input  [31:0] input_w,
    output [31:0] output_x
);

assign output_x = input_w;

endmodule